library ieee; --** allows use of the std_logic_vector type
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity g04_permutation is
port (input_code: in std_logic_vector(4 downto 0);
		rotor_type: in std_logic_vector(1 downto 0);
		output_code: out std_logic_vector(4 downto 0);
		inv_output_code: out std_logic_vector(4 downto 0));
end g04_permutation;
architecture behav of g04_permutation is
signal temp_inv_output_code, temp_output_code: std_logic_vector(4 downto 0);

begin
process(input_code,rotor_type)
begin
case rotor_type is
when "00" =>
	case input_code is
		when "00000"=>--**A**
			temp_output_code <= "00100";--**E**
			temp_inv_output_code <= "10100";--**U**
		when "00001"=>--**B**
			temp_output_code <= "01010";--**K**
			temp_inv_output_code <= "10110";--**W**
		when "00010"=>--**C**
			temp_output_code <= "01100";--**M**
			temp_inv_output_code <= "11000";--**Y**
		when "00011"=>--**D**
			temp_output_code <= "00101";--**F**
			temp_inv_output_code <= "00110";--**G**
		when "00100"=>--**E**
			temp_output_code <= "01011";--**L**
			temp_inv_output_code <= "00000";--**A**
		when "00101"=>--**F**
			temp_output_code <= "00110";--**G**
			temp_inv_output_code <= "00011";--**D**
		when "00110"=>--**G**
			temp_output_code <= "00011";--**D**
		   temp_inv_output_code <= "00101";--**F**
		when "00111"=>--**H**
			temp_output_code <= "10000";--**Q**
     		temp_inv_output_code <= "01111";--**P**
		when "01000"=>--**I**
			temp_output_code <= "10101";--**V**
			temp_inv_output_code <= "10101";--**V**
		when "01001"=>--**J**
			temp_output_code <= "11001";--**Z**
			temp_inv_output_code <= "11001";--**Z**
		when "01010"=>--**K**
			temp_output_code <= "01101";--**N**
			temp_inv_output_code <= "00001";--**B**
		when "01011"=>--**L**
			temp_output_code <= "10011";--**T**
			temp_inv_output_code <= "00100";--**E**
		when "01100"=>--**M**
			temp_output_code <= "01110";--**O**
			temp_inv_output_code <= "00010";--**C**
		when "01101"=>--**N**
			temp_output_code <= "10110"; --**W**
			temp_inv_output_code <= "01010";--**K**
		when "01110"=>--**O**
			temp_output_code <= "11000"; --**Y**
			temp_inv_output_code <= "01100";--**M**	
		when "01111"=>--**P**
			temp_output_code <= "00111"; --**H**
			temp_inv_output_code <= "10011";--**T**
		when "10000"=>--**Q**
			temp_output_code <= "10111"; --**X**
			temp_inv_output_code <= "00111";--**H**
		when "10001"=>--**R**
			temp_output_code <= "10100"; --**U**
			temp_inv_output_code <= "10111";--**X**					 
		when "10010"=>--**S**
			temp_output_code <= "10010"; --**S**
			temp_inv_output_code <= "10010";--**S**
		when "10011"=>--**T**
			temp_output_code <= "01111"; --**P**
			temp_inv_output_code <= "01011";--**L**	
		when "10100"=>--**U**
			temp_output_code <= "00000"; --**A**
			temp_inv_output_code <= "10001";--**R**
		when "10101"=>--**V**
			temp_output_code <= "01000"; --**I**
			temp_inv_output_code <= "01000";--**I**
		when "10110"=>--**W**
			temp_output_code <= "00001"; --**B**
			temp_inv_output_code <= "01101";--**N**		
		when "10111"=>--**X**
			temp_output_code <= "10001"; --**R**
			temp_inv_output_code <= "10000";--**Q**
		when "11000"=>--**Y**
			temp_output_code <= "00010"; --**C**
			temp_inv_output_code <= "01110";--**O**	
		when others=>--**Z**
			temp_output_code <= "01001"; --**J**
			temp_inv_output_code <= "01001";--**J**
END CASE;
when"01" =>			
	case input_code is
		when "00000"=>--**A**
			temp_output_code <= "00000";--**A**
			temp_inv_output_code <= "00000";--**A**
		when "00001"=>--**B**
			temp_output_code <= "01001";--**J**
			temp_inv_output_code <= "01001";--**J**
		when "00010"=>--**C**
			temp_output_code <= "00011";--**D**
			temp_inv_output_code <= "01111";--**P**
		when "00011"=>--**D**
			temp_output_code <= "01010";--**K**
			temp_inv_output_code <= "00010";--**C**
		when "00100"=>--**E**
			temp_output_code <= "10010";--**S**
			temp_inv_output_code <= "11001";--**Z**
		when "00101"=>--**F**
			temp_output_code <= "01000";--**I**
			temp_inv_output_code <= "10110";--**W**
		when "00110"=>--**G**
			temp_output_code <= "10001";--**R**
		   temp_inv_output_code <= "10001";--**R**
		when "00111"=>--**H**
			temp_output_code <= "10100";--**U**
     		temp_inv_output_code <= "01011";--**L**
		when "01000"=>--**I**
			temp_output_code <= "10111";--**X**
			temp_inv_output_code <= "00101";--**F**
		when "01001"=>--**J**
			temp_output_code <= "00001";--**B**
			temp_inv_output_code <= "00001";--**B**
		when "01010"=>--**K**
			temp_output_code <= "01011";--**L**
			temp_inv_output_code <= "00011";--**D**
		when "01011"=>--**L**
			temp_output_code <= "00111";--**H**
			temp_inv_output_code <= "01010";--**K**
		when "01100"=>--**M**
			temp_output_code <= "10110";--**W**
			temp_inv_output_code <= "01110";--**O**
		when "01101"=>--**N**
			temp_output_code <= "10011"; --**T**
			temp_inv_output_code <= "10011";--**T**
		when "01110"=>--**O**
			temp_output_code <= "01100"; --**M**
			temp_inv_output_code <= "11000";--**Y**	
		when "01111"=>--**P**
			temp_output_code <= "00010"; --**C**
			temp_inv_output_code <= "10100";--**U**
		when "10000"=>--**Q**
			temp_output_code <= "10000"; --**Q**
			temp_inv_output_code <= "10000";--**Q**
		when "10001"=>--**R**
			temp_output_code <= "00110"; --**G**
			temp_inv_output_code <= "00110";--**G**					 
		when "10010"=>--**S**
			temp_output_code <= "11001"; --**Z**
			temp_inv_output_code <= "00100";--**E**
		when "10011"=>--**T
			temp_output_code <= "01101"; --**N**
			temp_inv_output_code <= "01101";--**N**	
		when "10100"=>--**U**
			temp_output_code <= "01111"; --**P**
			temp_inv_output_code <= "00111";--**H**
		when "10101"=>--**V**
			temp_output_code <= "11000"; --**Y**
			temp_inv_output_code <= "10111";--**X**
		when "10110"=>--**W**
			temp_output_code <= "00101"; --**F**
			temp_inv_output_code <= "01100";--**M**		
		when "10111"=>--**X**
			temp_output_code <= "10101"; --**V**
			temp_inv_output_code <= "01000";--**I**
		when "11000"=>--**Y**
			temp_output_code <= "01110"; --**O**
			temp_inv_output_code <= "10101";--**V**	
		when others=>--**Z**
			temp_output_code <= "00100"; --**E**
			temp_inv_output_code <= "10010";--**S**
END CASE;
when"10" =>			
	case input_code is
		when "00000"=>--**A**
			temp_output_code <= "00001";--**B**
			temp_inv_output_code <= "10011";--**T**
		when "00001"=>--**B**
			temp_output_code <= "00011";--**D**
			temp_inv_output_code <= "00000";--**A**
		when "00010"=>--**C**
			temp_output_code <= "00101";--**F**
			temp_inv_output_code <= "00110";--**G**
		when "00011"=>--**D**
			temp_output_code <= "00111";--**H**
			temp_inv_output_code <= "00001";--**B**
		when "00100"=>--**E**
			temp_output_code <= "01001";--**J**
			temp_inv_output_code <= "01111";--**P**
		when "00101"=>--**F**
			temp_output_code <= "01011";--**L**
			temp_inv_output_code <= "00010";--**C**
		when "00110"=>--**G**
			temp_output_code <= "00010";--**C**
		   temp_inv_output_code <= "10010";--**S**
		when "00111"=>--**H**
			temp_output_code <= "01111";--**P**
     		temp_inv_output_code <= "00011";--**D**
		when "01000"=>--**I**
			temp_output_code <= "10001";--**R**
			temp_inv_output_code <= "10000";--**Q**
		when "01001"=>--**J**
			temp_output_code <= "10011";--**T**
			temp_inv_output_code <= "00100";--**E**
		when "01010"=>--**K**
			temp_output_code <= "10111";--**X**
			temp_inv_output_code <= "10100";--**U**
		when "01011"=>--**L**
			temp_output_code <= "10101";--**V**
			temp_inv_output_code <= "00101";--**F**
		when "01100"=>--**M**
			temp_output_code <= "11001";--**Z**
			temp_inv_output_code <= "10101";--**V**
		when "01101"=>--**N**
			temp_output_code <= "01101"; --**N**
			temp_inv_output_code <= "01101";--**N**
		when "01110"=>--**O**
			temp_output_code <= "11000"; --**Y**
			temp_inv_output_code <= "11001";--**Z**	
		when "01111"=>--**P**
			temp_output_code <= "00100"; --**E**
			temp_inv_output_code <= "00111";--**H**
		when "10000"=>--**Q**
			temp_output_code <= "01000"; --**I**
			temp_inv_output_code <= "11000";--**Y**
		when "10001"=>--**R**
			temp_output_code <= "10110"; --**W**
			temp_inv_output_code <= "01000";--**I**					 
		when "10010"=>--**S**
			temp_output_code <= "00110"; --**G**
			temp_inv_output_code <= "10111";--**X**
		when "10011"=>--**T
			temp_output_code <= "00000"; --**A**
			temp_inv_output_code <= "01010";--**J**	
		when "10100"=>--**U**
			temp_output_code <= "01010"; --**K**
			temp_inv_output_code <= "10110";--**W**
		when "10101"=>--**V**
			temp_output_code <= "01100"; --**M**
			temp_inv_output_code <= "01011";--**L**
		when "10110"=>--**W**
			temp_output_code <= "10100"; --**U**
			temp_inv_output_code <= "10001";--**R**		
		when "10111"=>--**X**
			temp_output_code <= "10001"; --**S**
			temp_inv_output_code <= "01010";--**K**
		when "11000"=>--**Y**
			temp_output_code <= "10000"; --**Q**
			temp_inv_output_code <= "01110";--**O**	
		when others=>--**Z**
			temp_output_code <= "01110"; --**O**
			temp_inv_output_code <= "01100";--**M**
END CASE;
when others =>			
	case input_code is
		when "00000"=>--**A**
			temp_output_code <= "00100";--**E**
			temp_inv_output_code <= "00111";--**H**
		when "00001"=>--**B**
			temp_output_code <= "10010";--**S**
			temp_inv_output_code <= "11001";--**Z**
		when "00010"=>--**C**
			temp_output_code <= "01110";--**O**
			temp_inv_output_code <= "10110";--**W**
		when "00011"=>--**D**
			temp_output_code <= "10101";--**V**
			temp_inv_output_code <= "10101";--**V**
		when "00100"=>--**E**
			temp_output_code <= "01111";--**P**
			temp_inv_output_code <= "00000";--**A**
		when "00101"=>--**F**
			temp_output_code <= "11001";--**Z**
			temp_inv_output_code <= "10001";--**R**
		when "00110"=>--**G**
			temp_output_code <= "01001";--**J**
		   temp_inv_output_code <= "10011";--**T**
		when "00111"=>--**H**
			temp_output_code <= "00000";--**A**
     		temp_inv_output_code <= "01101";--**N**
		when "01000"=>--**I**
			temp_output_code <= "11000";--**Y**
			temp_inv_output_code <= "01011";--**L**
		when "01001"=>--**J**
			temp_output_code <= "10000";--**Q**
			temp_inv_output_code <= "00110";--**G**
		when "01010"=>--**K**
			temp_output_code <= "10100";--**U**
			temp_inv_output_code <= "10100";--**U**
		when "01011"=>--**L**
			temp_output_code <= "01000";--**I**
			temp_inv_output_code <= "01111";--**P**
		when "01100"=>--**M**
			temp_output_code <= "10001";--**R**
			temp_inv_output_code <= "10111";--**X**
		when "01101"=>--**N**
			temp_output_code <= "00111"; --**H**
			temp_inv_output_code <= "10000";--**Q**
		when "01110"=>--**O**
			temp_output_code <= "10111"; --**X**
			temp_inv_output_code <= "00010";--**C**	
		when "01111"=>--**P**
			temp_output_code <= "01011"; --**L**
			temp_inv_output_code <= "00100";--**E**
		when "10000"=>--**Q**
			temp_output_code <= "01101"; --**N**
			temp_inv_output_code <= "01001";--**J**
		when "10001"=>--**R**
			temp_output_code <= "00101"; --**F**
			temp_inv_output_code <= "01100";--**M**					 
		when "10010"=>--**S**
			temp_output_code <= "10011"; --**T**
			temp_inv_output_code <= "00001";--**B**
		when "10011"=>--**T
			temp_output_code <= "00110"; --**G**
			temp_inv_output_code <= "10010";--**S**	
		when "10100"=>--**U**
			temp_output_code <= "01010"; --**K**
			temp_inv_output_code <= "01010";--**K**
		when "10101"=>--**V**
			temp_output_code <= "00011"; --**D**
			temp_inv_output_code <= "00011";--**D**
		when "10110"=>--**W**
			temp_output_code <= "00010"; --**C**
			temp_inv_output_code <= "11000";--**Y**		
		when "10111"=>--**X**
			temp_output_code <= "01100"; --**M**
			temp_inv_output_code <= "01110";--**0**
		when "11000"=>--**Y**
			temp_output_code <= "10110"; --**W**
			temp_inv_output_code <= "01000";--**I**	
		when others=>--**Z**
			temp_output_code <= "00001"; --**B**
			temp_inv_output_code <= "00101";--**F**
END CASE;
END CASE;
END PROCESS;
output_code<= temp_output_code;
inv_output_code<= temp_inv_output_code;
END behav;
